module constantvaluegenerator_project(output wire[width-1:0] databus);

	parameter width=4;
	parameter value=1;
	assign databus = 4;
	
endmodule